`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01.08.2025 18:10:52
// Design Name: 
// Module Name: aes
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module aes(clk, reset, in, key, ciphertext);
    input logic clk, reset;
    input logic [127:0] in;
    input logic [127:0] key;
    output logic [127:0] ciphertext;
    
    logic [7:0] keyMatrix [0:3][0:3];
    logic [7:0] inputBlock [0:3][0:3];

    
    // states after each round
    logic [7:0] state0      [0:3][0:3];
    logic [7:0] state1      [0:3][0:3];
    logic [7:0] state2      [0:3][0:3];
    logic [7:0] state3      [0:3][0:3];
    logic [7:0] state4      [0:3][0:3];
    logic [7:0] state5      [0:3][0:3];
    logic [7:0] state6      [0:3][0:3];
    logic [7:0] state7      [0:3][0:3];
    logic [7:0] state8      [0:3][0:3];
    logic [7:0] state9      [0:3][0:3];
    logic [7:0] state10      [0:3][0:3];
    
    // temp vars to store states
    logic [7:0] op1_out      [0:3][0:3];
    logic [7:0] op2_out      [0:3][0:3];
    logic [7:0] op3_out      [0:3][0:3];
    logic [7:0] op4_out      [0:3][0:3];
    logic [7:0] op5_out      [0:3][0:3];
    logic [7:0] op6_out      [0:3][0:3];
    logic [7:0] op7_out      [0:3][0:3];
    logic [7:0] op8_out      [0:3][0:3];
    logic [7:0] op9_out      [0:3][0:3];
    logic [7:0] op10_out      [0:3][0:3];
    
    // keys generated by key Expansion module
    
    logic [7:0] key0      [0:3][0:3];
    logic [7:0] key1      [0:3][0:3];
    logic [7:0] key2      [0:3][0:3];
    logic [7:0] key3      [0:3][0:3];
    logic [7:0] key4      [0:3][0:3];
    logic [7:0] key5      [0:3][0:3];
    logic [7:0] key6      [0:3][0:3];
    logic [7:0] key7      [0:3][0:3];
    logic [7:0] key8      [0:3][0:3];
    logic [7:0] key9      [0:3][0:3];
    logic [7:0] key10      [0:3][0:3];

    
    
    keyExpander KeyExpansion(.key(key), .key0(key0), .key1(key1), .key2(key2), .key3(key3), .key4(key4), .key5(key5), .key6(key6), .key7(key7), .key8(key8), .key9(key9), .key10(key10));
    
    operations op1(.in(state0), .key(key1), .out(op1_out));
    operations op2(.in(state1), .key(key2), .out(op2_out));
    operations op3(.in(state2), .key(key3), .out(op3_out));
    operations op4(.in(state3), .key(key4), .out(op4_out));
    operations op5(.in(state4), .key(key5), .out(op5_out));
    operations op6(.in(state5), .key(key6), .out(op6_out));
    operations op7(.in(state6), .key(key7), .out(op7_out));
    operations op8(.in(state7), .key(key8), .out(op8_out));
    operations op9(.in(state8), .key(key9), .out(op9_out));
    operationN op10(.in(state9), .key(key10), .out(op10_out));
    
    
    always_ff @(posedge clk or posedge reset) begin 
        if(reset) begin        
            for (int j = 0; j < 4; j++) begin  
                for (int i = 0; i < 4; i++) begin 
                    inputBlock[i][j] = in[127 - ((4 * j + i) * 8) -: 8];
                end
            end
        end
    end
       
   
    always_ff @(posedge clk or posedge reset) begin // ROUND 0
        if(!reset) begin
            foreach (state0[i,j])
               state0[i][j] <= key0[i][j] ^ inputBlock[i][j];

        end
    end
    
    always_ff @(posedge clk or posedge reset) begin // ROUND 1
        if(!reset) begin
            foreach (state1[i,j])
               state1[i][j] <= op1_out[i][j];
        end
    end
    
    always_ff @(posedge clk or posedge reset) begin // ROUND 2
        if(!reset) begin
            foreach (state2[i,j])
               state2[i][j] <= op2_out[i][j];
        end
    end
    
    
    always_ff @(posedge clk or posedge reset) begin // ROUND 3
        if(!reset) begin
            foreach (state3[i,j])
               state3[i][j] <= op3_out[i][j];
        end
    end
    
    
    always_ff @(posedge clk or posedge reset) begin // ROUND 4
        if(!reset) begin
            foreach (state4[i,j])
               state4[i][j] <= op4_out[i][j];
        end
    end
    
    
    always_ff @(posedge clk or posedge reset) begin // ROUND 5
        if(!reset) begin
            foreach (state5[i,j])
               state5[i][j] <= op5_out[i][j];
        end
    end
    
    
    always_ff @(posedge clk or posedge reset) begin // ROUND 6
        if(!reset) begin
            foreach (state6[i,j])
               state6[i][j] <= op6_out[i][j];
        end
    end
    
    
    always_ff @(posedge clk or posedge reset) begin // ROUND 7
        if(!reset) begin
            foreach (state7[i,j])
               state7[i][j] <= op7_out[i][j];
        end
    end
    
    always_ff @(posedge clk or posedge reset) begin // ROUND 8
        if(!reset) begin
            foreach (state8[i,j])
               state8[i][j] <= op8_out[i][j];
        end
    end
    
    always_ff @(posedge clk or posedge reset) begin // ROUND 9
        if(!reset) begin
            foreach (state9[i,j])
               state9[i][j] <= op9_out[i][j];
        end
    end
    
    always_ff @(posedge clk or posedge reset) begin // ROUND 10
        if(!reset) begin
            foreach (state10[i,j])
               state10[i][j] <= op10_out[i][j];
               
            for (int k = 0; k < 4; k++) begin
                for (int m = 0; m < 4; m++) begin
                    ciphertext[127 - ((4*k + m)*8) -: 8] <= op10_out[m][k];
                end
            end
        end
    end

endmodule
